--
-- Equality comparator template.
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Buf_7 is
  generic(BusWidth : integer := 7);
  port(
        --Data signals.
        i : in std_logic_vector(BusWidth - 1 downto 0);
        o : out std_logic_vector(BusWidth - 1 downto 0)
      );
end Buf_7;

architecture Behavioral of Buf_7 is
begin
  o <= i;
end Behavioral;

